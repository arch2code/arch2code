//copyright Arch2Code authors 2024

// GENERATED_CODE_PARAM --block=simple --parentModule
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
// GENERATED_CODE_END
