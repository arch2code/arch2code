// GENERATED_CODE_PARAM --block=blockBX
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
//module as defined by block: blockBX
module blockBX
// Generated Import package statement(s)
import hierInclude_package::*;
import hierIncludeB_package::*;
(
    rdy_vld_if.src bx2y,
    rdy_vld_if.src bx2z,
    rdy_vld_if.dst anInterface,
    req_ack_if.src b2C,
    input clk, rst_n
);

    // Interface Instances, needed for between instanced modules inside this module

// Instances

// GENERATED_CODE_END

endmodule: blockBX