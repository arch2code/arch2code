// GENERATED_CODE_PARAM --block=blockD
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
//module as defined by block: blockD
module blockD
// Generated Import package statement(s)
import mixedInclude_package::*;
import mixedBlockC_package::*;
import mixed_package::*;
(
    rdy_vld_if.src cStuffIf,
    rdy_vld_if.src dee0,
    rdy_vld_if.src dee1,
    rdy_vld_if.src outD,
    rdy_vld_if.dst inD,
    req_ack_if.dst btod,
    status_if.dst rwD,
    status_if.src roBsize,
    memory_if.src blockBTable1,
    memory_if.src blockBTableSP,
    input clk, rst_n
);

    // Interface Instances, needed for between instanced modules inside this module

// Instances
// GENERATED_CODE_END

endmodule: blockD
