`ifndef _PIPE_HDL_SV_WRAPPER_SV_GUARD_
`define _PIPE_HDL_SV_WRAPPER_SV_GUARD_

// GENERATED_CODE_PARAM --block=pipe
// GENERATED_CODE_BEGIN --template=module_hdl_sv_wrapper
// GENERATED_CODE_END

`endif // _PIPE_HDL_SV_WRAPPER_SV_GUARD_
