// GENERATED_CODE_PARAM --block=cpu
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
//module as defined by block: cpu
module cpu
// Generated Import package statement(s)
import mixed_package::*;
(
    apb_if.src apbReg,
    input clk, rst_n
);

    // Interface Instances, needed for between instanced modules inside this module


// Instances
// GENERATED_CODE_END

endmodule: cpu