// GENERATED_CODE_PARAM --block=inAndOut
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
//module as defined by block: inAndOut
module inAndOut
// Generated Import package statement(s)
import inAndOut_package::*;
(
    rdy_vld_if.src aOut,
    rdy_vld_if.dst aIn,
    req_ack_if.src bOut,
    req_ack_if.dst bIn,
    pop_ack_if.src dOut,
    pop_ack_if.dst dIn,
    input clk, rst_n
);

    // Interface Instances, needed for between instanced modules inside this module


// Instances
// GENERATED_CODE_END

endmodule: inAndOut