// GENERATED_CODE_PARAM --contexts hierIncludeNestedTop.yaml
// GENERATED_CODE_BEGIN --template=package --fileMapKey=package_sv
package hierIncludeNestedTop_package;
//constants as defined by the scope of the following context(s): ('hierIncludeNestedTop.yaml',)
//         YET_ANOTHER_SIZE =                   'd8;  // The size of yet another size
localparam YET_ANOTHER_SIZE =                 32'h0000_0008;  // The size of yet another size

// types

// enums

// structures
endpackage : hierIncludeNestedTop_package
// GENERATED_CODE_END
