// GENERATED_CODE_PARAM --context mixedInclude.yaml
// GENERATED_CODE_BEGIN --template=package --fileMapKey=package_sv
package mixedInclude_package;
// Generated Import package statement(s)
import mixedNestedInclude_package::*;
localparam int unsigned BSIZE = 32'h0000_000A;  // The size of B, used for memory wordlines
localparam int unsigned BSIZE_LOG2 = 32'h0000_0004;  // The size of B, used for memory wordlines log 2

// types

// enums

// structures
endpackage : mixedInclude_package
// GENERATED_CODE_END
