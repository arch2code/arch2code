// GENERATED_CODE_PARAM --block=consumer
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
//module as defined by block: consumer
module consumer
// Generated Import package statement(s)
import axiDemo_package::*;
(
    axi_read_if.dst axiRd0,
    axi_read_if.dst axiRd1,
    axi_read_if.dst axiRd2,
    axi_read_if.dst axiRd3,
    axi_write_if.dst axiWr0,
    axi_write_if.dst axiWr1,
    axi_write_if.dst axiWr2,
    axi_write_if.dst axiWr3,
    axi4_stream_if.dst axiStr0,
    axi4_stream_if.dst axiStr1,
    input clk, rst_n
);

    // Interface Instances, needed for between instanced modules inside this module

// Instances

// GENERATED_CODE_END

endmodule: consumer
