../../../../../../../examples/axiDemo/systemVerilog/producer.sv