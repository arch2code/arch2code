../../../../../../../examples/axiDemo/systemVerilog/top.sv