../../../../../../../examples/axiDemo/systemVerilog/consumer.sv