// GENERATED_CODE_PARAM --context b/hierIncludeBInclude.yaml
// GENERATED_CODE_BEGIN --template=package --fileMapKey=package_sv
package hierIncludeBInclude_package;
localparam int B_ANOTHER_SIZE = 32'h0000_0009;  // The size for b another size

// types

// enums

// structures
endpackage : hierIncludeBInclude_package
// GENERATED_CODE_END
