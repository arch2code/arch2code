
// copyright Arch2Code authors 2024
// GENERATED_CODE_PARAM --contexts=simple/simple.yaml
// GENERATED_CODE_BEGIN --template=package --fileMapKey=package_sv
// GENERATED_CODE_END
