// GENERATED_CODE_PARAM --contexts b/hierIncludeBInclude.yaml
// GENERATED_CODE_BEGIN --template=package --fileMapKey=package_sv
package hierIncludeBInclude_package;
//constants as defined by the scope of the following context(s): ('b/hierIncludeBInclude.yaml',)
//         B_ANOTHER_SIZE =                     'd9;  // The size for b another size
localparam B_ANOTHER_SIZE =                   32'h0000_0009;  // The size for b another size

// types

// enums

// structures
endpackage : hierIncludeBInclude_package
// GENERATED_CODE_END
