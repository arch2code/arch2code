`ifndef _SIMPLE_HDL_SV_WRAPPER_SV_GUARD_
`define _SIMPLE_HDL_SV_WRAPPER_SV_GUARD_

// GENERATED_CODE_PARAM --block=simple
// GENERATED_CODE_BEGIN --template=module_hdl_sv_wrapper
// GENERATED_CODE_END

`endif // _SIMPLE_HDL_SV_WRAPPER_SV_GUARD_
