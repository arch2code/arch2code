// GENERATED_CODE_PARAM --context hierIncludeTop.yaml
// GENERATED_CODE_BEGIN --template=package --fileMapKey=package_sv
package hierIncludeTop_package;
// Generated Import package statement(s)
import hierIncludeNestedTop_package::*;
localparam int unsigned ANOTHER_SIZE = 32'h0000_0004;  // The size for another size

// types

// enums

// structures
endpackage : hierIncludeTop_package
// GENERATED_CODE_END
