// GENERATED_CODE_PARAM --context c/hierIncludeC.yaml
// GENERATED_CODE_BEGIN --template=package --fileMapKey=package_sv
package hierIncludeC_package;
// Generated Import package statement(s)
import hierIncludeTop_package::*;
import hierInclude_package::*;
import hierIncludeCInclude_package::*;

// types
typedef logic[C_ANOTHER_SIZE-1:0] cSizeT; //A type from an include

// enums

// structures
typedef struct packed {
    cSizeT cAnother; //
} cSt;

endpackage : hierIncludeC_package
// GENERATED_CODE_END
