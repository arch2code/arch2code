// GENERATED_CODE_PARAM --block=cpu --parentModule
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
//module as defined by block: cpu
module cpu
// Generated Import package statement(s)
import apbDecode_package::*;
(
    apb_if.src apbReg,
    input clk, rst_n
);

    // Interface Instances, needed for between instanced modules inside this module

// Instances
endmodule // cpu
// GENERATED_CODE_END
