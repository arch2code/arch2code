// GENERATED_CODE_PARAM --context mixedNestedInclude.yaml
// GENERATED_CODE_BEGIN --template=package --fileMapKey=package_sv
package mixedNestedInclude_package;
//         DSIZE =                              'd1;  // The size of D
localparam DSIZE =                            32'h0000_0001;  // The size of D
//         DSIZE2 =                             'd2;  // The size of D2
localparam DSIZE2 =                           32'h0000_0002;  // The size of D2

// types

// enums

// structures
endpackage : mixedNestedInclude_package
// GENERATED_CODE_END
