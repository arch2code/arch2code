../../../../../../examples/mixed/systemVerilog/blockB.sv