`ifndef VL_WRAP_SV_
`define VL_WRAP_SV_

`include "blockA_hdl_sv_wrapper.sv"
`include "blockF_uBlockF0_hdl_sv_wrapper.sv"
`include "blockF_uBlockF1_hdl_sv_wrapper.sv"

`endif // VL_WRAP_SV_
