// GENERATED_CODE_PARAM --block=blockBY --parentModule
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
//module as defined by block: blockBY
module blockBY
// Generated Import package statement(s)
import hierIncludeB_package::*;
(
    rdy_vld_if.dst x,
    input clk, rst_n
);

    // Interface Instances, needed for between instanced modules inside this module

// Instances
endmodule // blockBY
// GENERATED_CODE_END
