`ifndef VL_WRAP_SV_
`define VL_WRAP_SV_

`include "blockA_hdl_sv_wrapper.sv"
`include "blockB_hdl_sv_wrapper.sv"
`include "apbDecode_hdl_sv_wrapper.sv"
`include "someRapper_hdl_sv_wrapper.sv"

`endif // VL_WRAP_SV_
