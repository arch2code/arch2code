// GENERATED_CODE_PARAM --block=blockA
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
//module as defined by block: blockA
module blockA
// Generated Import package statement(s)
import hierInclude_package::*;
(
    rdy_vld_if.src anInterfaceB,
    rdy_vld_if.src anInterfaceC,
    input clk, rst_n
);

    // Interface Instances, needed for between instanced modules inside this module


// Instances
// GENERATED_CODE_END

endmodule: blockA