`ifndef VL_WRAP_SV_
`define VL_WRAP_SV_

`include "producer_hdl_sv_wrapper.sv"
`include "consumer_hdl_sv_wrapper.sv"

`endif // VL_WRAP_SV_
