// GENERATED_CODE_PARAM --block=blockC
// GENERATED_CODE_BEGIN --template=moduleInterfacesInstances
//module as defined by block: blockC
module blockC
// Generated Import package statement(s)
import mixedBlockC_package::*;
(
    rdy_vld_if.dst see,
    input clk, rst_n
);

    // Interface Instances, needed for between instanced modules inside this module

// Instances

// GENERATED_CODE_END

endmodule: blockC

